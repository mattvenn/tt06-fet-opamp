* NGSPICE file created from opamp_parax.ext - technology: sky130A

.subckt opamp_parax VDD ZREF vin_n vin_p Vout VGND
R0 ZREF VGND sky130_fd_pr__res_generic_l1 w=1 l=5
X0 a_n874_n1404# a_n874_n1404# VGND.t6 VGND.t5 sky130_fd_pr__nfet_01v8 ad=1.74 pd=12.58 as=0 ps=0 w=6 l=0.6
**devattr s=69600,2516 d=69600,2516
X1 Vout.t1 a_728_n1284# VGND.t2 VGND.t1 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=6 l=0.6
**devattr s=69600,2516 d=69600,2516
X2 VDD.t5 VGND.t7 w_n1008_n1084# VDD.t4 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=1.74 ps=12.58 w=6 l=0.6
**devattr s=69600,2516 d=69600,2516
X3 w_n1008_n1084# vin_p.t0 a_728_n1284# w_n1008_n1084# sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=0.6
**devattr s=69600,2516 d=69600,2516
X4 a_2502_n1184.t1 Vout.t0 sky130_fd_pr__cap_mim_m3_1 l=15 w=17.55
X5 VDD.t3 VGND.t8 Vout.t2 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=6 l=0.6
**devattr s=69600,2516 d=69600,2516
X6 VDD.t1 VGND.t9 ZREF.t0 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=6 l=0.6
**devattr s=69600,2516 d=69600,2516
X7 a_728_n1284# a_n874_n1404# VGND.t4 VGND.t3 sky130_fd_pr__nfet_01v8 ad=1.74 pd=12.994286 as=0 ps=0 w=6 l=0.6
**devattr s=69600,2516 d=69600,2516
X8 a_2502_n1184.t0 VDD.t6 a_728_n1284# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.29 ps=2.165714 w=1 l=0.6
**devattr s=11600,516 d=11600,516
R1 VDD ZREF sky130_fd_pr__res_generic_l1 w=1 l=5
X9 w_n1008_n1084# vin_n.t0 a_n874_n1404# w_n1008_n1084# sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=0.6
**devattr s=69600,2516 d=69600,2516
R2 VGND.n49 VGND.n48 31557.4
R3 VGND.n38 VGND.n34 17132.9
R4 VGND.n33 VGND.n30 5463.85
R5 VGND.n40 VGND.n30 5463.85
R6 VGND.n33 VGND.n31 5463.85
R7 VGND.n40 VGND.n31 5463.85
R8 VGND.n21 VGND.n7 5463.85
R9 VGND.n50 VGND.n5 5463.85
R10 VGND.n50 VGND.n6 5463.85
R11 VGND.n21 VGND.n8 5463.85
R12 VGND.n11 VGND.n7 4386.15
R13 VGND.n11 VGND.n5 4386.15
R14 VGND.n12 VGND.n8 4386.15
R15 VGND.n12 VGND.n6 4386.15
R16 VGND.n36 VGND.n24 2566.79
R17 VGND.n47 VGND.n24 2566.79
R18 VGND.n36 VGND.n25 2566.79
R19 VGND.n47 VGND.n25 2566.79
R20 VGND.n14 VGND.n11 1077.71
R21 VGND.n14 VGND.n12 1077.71
R22 VGND.n22 VGND.t3 784.087
R23 VGND.n13 VGND.t3 784.087
R24 VGND.n13 VGND.t5 784.087
R25 VGND.n49 VGND.t5 784.087
R26 VGND.n34 VGND.t1 679.755
R27 VGND.n39 VGND.t1 679.755
R28 VGND.n48 VGND.n23 488.599
R29 VGND.n32 VGND.n29 355.012
R30 VGND.n41 VGND.n29 355.012
R31 VGND.n32 VGND.n28 355.012
R32 VGND.n20 VGND.n9 355.012
R33 VGND.n51 VGND.n4 355.012
R34 VGND.n23 VGND.n22 353.202
R35 VGND.n52 VGND.n51 349.365
R36 VGND.n42 VGND.n41 347.483
R37 VGND.n20 VGND.n19 344.848
R38 VGND.n10 VGND.n9 284.988
R39 VGND.n10 VGND.n4 284.988
R40 VGND.n17 VGND.n16 284.988
R41 VGND.n16 VGND.n3 284.988
R42 VGND.n0 VGND.t8 228.256
R43 VGND.n0 VGND.t7 213.042
R44 VGND.n1 VGND.t9 213.042
R45 VGND.n37 VGND.n36 185.922
R46 VGND.n35 VGND.n26 166.776
R47 VGND.n35 VGND.n27 166.776
R48 VGND.n46 VGND.n26 166.776
R49 VGND.n46 VGND.n45 166.4
R50 VGND.n37 VGND.t0 150.575
R51 VGND.n41 VGND.n40 146.25
R52 VGND.n40 VGND.n39 146.25
R53 VGND.n33 VGND.n32 146.25
R54 VGND.n34 VGND.n33 146.25
R55 VGND.n26 VGND.n24 146.25
R56 VGND.t0 VGND.n24 146.25
R57 VGND.n27 VGND.n25 146.25
R58 VGND.t0 VGND.n25 146.25
R59 VGND.n15 VGND.n14 146.25
R60 VGND.n14 VGND.n13 146.25
R61 VGND.n21 VGND.n20 146.25
R62 VGND.n22 VGND.n21 146.25
R63 VGND.n51 VGND.n50 146.25
R64 VGND.n50 VGND.n49 146.25
R65 VGND.n47 VGND.n46 117.001
R66 VGND.n48 VGND.n47 117.001
R67 VGND.n36 VGND.n35 117.001
R68 VGND.n15 VGND.n10 70.024
R69 VGND.n16 VGND.n15 70.024
R70 VGND.n39 VGND.n38 47.5923
R71 VGND.n38 VGND.n37 33.3793
R72 VGND.n31 VGND.n28 29.2505
R73 VGND.t1 VGND.n31 29.2505
R74 VGND.n30 VGND.n29 29.2505
R75 VGND.t1 VGND.n30 29.2505
R76 VGND.n9 VGND.n7 29.2505
R77 VGND.n7 VGND.t3 29.2505
R78 VGND.n5 VGND.n4 29.2505
R79 VGND.t5 VGND.n5 29.2505
R80 VGND.n6 VGND.n3 29.2505
R81 VGND.t5 VGND.n6 29.2505
R82 VGND.n17 VGND.n8 29.2505
R83 VGND.n8 VGND.t3 29.2505
R84 VGND.n55 VGND.n1 15.1666
R85 VGND.n18 VGND.t4 14.4211
R86 VGND.n53 VGND.t6 14.3926
R87 VGND.n43 VGND.t2 14.3699
R88 VGND.t0 VGND.n23 11.8683
R89 VGND.n19 VGND.n17 10.1652
R90 VGND.n45 VGND.n44 10.0105
R91 VGND.n42 VGND.n28 7.52991
R92 VGND.n52 VGND.n3 5.64756
R93 VGND.n44 VGND.n43 5.26544
R94 VGND.n1 VGND.n0 4.37237
R95 VGND.n19 VGND.n18 3.1005
R96 VGND.n54 VGND.n2 2.5824
R97 VGND.n53 VGND.n52 2.3255
R98 VGND.n44 VGND.n2 1.94544
R99 VGND.n43 VGND.n42 1.32907
R100 VGND.n55 VGND.n54 1.21171
R101 VGND.n45 VGND.n27 0.376971
R102 VGND VGND.n55 0.302375
R103 VGND.n18 VGND.n2 0.2615
R104 VGND.n54 VGND.n53 0.131
R105 Vout.n0 Vout.t2 39.9369
R106 Vout.n0 Vout.t1 14.5696
R107 Vout.n1 Vout.t0 2.58415
R108 Vout.n1 Vout.n0 1.39782
R109 Vout Vout.n1 0.336304
R110 VDD.n32 VDD.n5 3360
R111 VDD.n36 VDD.n3 3360
R112 VDD.n21 VDD.n15 3360
R113 VDD.n19 VDD.n18 3360
R114 VDD.n30 VDD.n8 2703.53
R115 VDD.n8 VDD.n3 2703.53
R116 VDD.n33 VDD.n32 2703.53
R117 VDD.n34 VDD.n33 2703.53
R118 VDD.t4 VDD.n7 1421.29
R119 VDD.n7 VDD.t0 1421.29
R120 VDD.n31 VDD.n5 1019.46
R121 VDD.n36 VDD.n35 1019.46
R122 VDD.n18 VDD.n17 1019.46
R123 VDD.n21 VDD.n20 1019.46
R124 VDD.n8 VDD.n4 656.471
R125 VDD.n33 VDD.n4 656.471
R126 VDD.n37 VDD.n2 358.401
R127 VDD.n9 VDD.n6 358.401
R128 VDD.n29 VDD.n9 358.401
R129 VDD.n22 VDD.n14 358.401
R130 VDD.n16 VDD.n14 358.401
R131 VDD.n16 VDD.n13 358.401
R132 VDD.n23 VDD.n22 350.495
R133 VDD.n38 VDD.n37 348.236
R134 VDD.n10 VDD.n6 288.377
R135 VDD.n10 VDD.n2 288.377
R136 VDD.n12 VDD.n1 288.377
R137 VDD.n28 VDD.n12 282.353
R138 VDD.n25 VDD.t6 114.528
R139 VDD.n12 VDD.n11 70.024
R140 VDD.n11 VDD.n10 70.024
R141 VDD.n11 VDD.n4 46.2505
R142 VDD.n7 VDD.n4 46.2505
R143 VDD.n37 VDD.n36 46.2505
R144 VDD.n9 VDD.n5 46.2505
R145 VDD.n22 VDD.n21 46.2505
R146 VDD.n18 VDD.n16 46.2505
R147 VDD.n24 VDD.t3 39.7606
R148 VDD.n0 VDD.t1 39.7543
R149 VDD.n26 VDD.t5 39.7543
R150 VDD.n38 VDD.n1 10.1652
R151 VDD.n34 VDD.n2 9.2505
R152 VDD.n32 VDD.n6 9.2505
R153 VDD.n32 VDD.t4 9.2505
R154 VDD.n30 VDD.n29 9.2505
R155 VDD.n3 VDD.n1 9.2505
R156 VDD.t0 VDD.n3 9.2505
R157 VDD.n19 VDD.n14 9.2505
R158 VDD.n15 VDD.n13 9.2505
R159 VDD.n23 VDD.n13 7.90638
R160 VDD.n31 VDD.n30 6.42675
R161 VDD.n35 VDD.n34 6.42675
R162 VDD.n17 VDD.n15 6.42675
R163 VDD.n20 VDD.n19 6.42675
R164 VDD.n29 VDD.n28 6.02403
R165 VDD.n35 VDD.t0 2.80756
R166 VDD.t4 VDD.n31 2.80756
R167 VDD.n20 VDD.t2 2.80756
R168 VDD.n17 VDD.t2 2.80756
R169 VDD.n28 VDD.n27 1.8605
R170 VDD.n25 VDD.n24 1.78992
R171 VDD.n39 VDD.n38 1.5505
R172 VDD.n24 VDD.n23 1.32907
R173 VDD.n26 VDD.n25 1.22396
R174 VDD.n27 VDD.n0 0.988864
R175 VDD VDD.n39 0.673909
R176 VDD.n39 VDD.n0 0.0120582
R177 VDD.n27 VDD.n26 0.00734932
R178 vin_p vin_p.t0 230.714
R179 a_2502_n1184.t0 a_2502_n1184.t1 89.7326
R180 ZREF ZREF.t0 131.24
R181 vin_n vin_n.t0 216.827
C0 vin_n vin_p 0.210606f
C1 li_n1228_n2039# w_n1008_n1084# 0.009085f
C2 a_n874_n1404# li_n1228_n981# 0.001658f
C3 li_n1228_n981# ZREF 0.179596f
C4 li_n1228_n2039# vin_n 0.014753f
C5 a_728_n1284# a_n874_n1404# 0.658987f
C6 w_n1008_n1084# li_n1228_n981# 0.129668f
C7 Vout a_728_n1284# 0.673923f
C8 vin_p li_n1228_n981# 0.151835f
C9 a_728_n1284# w_n1008_n1084# 0.759205f
C10 vin_n li_n1228_n981# 0.148464f
C11 VDD a_n874_n1404# 1.69e-19
C12 a_728_n1284# vin_p 0.642694f
C13 VDD ZREF 0.637682f
C14 VDD Vout 0.718665f
C15 VDD w_n1008_n1084# 0.911518f
C16 VDD vin_p 0.256783f
C17 VDD vin_n 0.002184f
C18 a_n874_n1404# ZREF 0.01426f
C19 Vout a_n874_n1404# 0.037248f
C20 w_n1008_n1084# a_n874_n1404# 0.736604f
C21 w_n1008_n1084# ZREF 0.026287f
C22 Vout w_n1008_n1084# 0.02174f
C23 VDD li_n1228_n981# 0.114337f
C24 vin_p a_n874_n1404# 0.018769f
C25 vin_n a_n874_n1404# 0.728268f
C26 vin_p ZREF 0.560099f
C27 Vout vin_p 0.00955f
C28 VDD a_728_n1284# 0.137643f
C29 vin_n ZREF 0.264221f
C30 Vout vin_n 0.004564f
C31 vin_p w_n1008_n1084# 1.93714f
C32 vin_n w_n1008_n1084# 1.08259f
C33 li_n1228_n2039# a_n874_n1404# 0.011878f
C34 li_n1228_n2039# ZREF 0.041726f
C35 vin_p VGND 1.20316f
C36 vin_n VGND 0.614746f
C37 Vout VGND 12.693263f
C38 ZREF VGND 2.38618f
C39 VDD VGND 15.896199f
C40 li_n1228_n2039# VGND 0.752214f $ **FLOATING
C41 li_n1228_n981# VGND 0.520365f $ **FLOATING
C42 a_728_n1284# VGND 2.90416f
C43 a_n874_n1404# VGND 3.17294f
C44 w_n1008_n1084# VGND 7.56163f
C45 a_2502_n1184.t1 VGND 24.4733f
C46 a_2502_n1184.t0 VGND 0.026705f
C47 Vout.t2 VGND 0.110597f
C48 Vout.t1 VGND 0.10775f
C49 Vout.n0 VGND 1.04598f
C50 Vout.t0 VGND 22.196001f
C51 Vout.n1 VGND 0.961303f
.ends

