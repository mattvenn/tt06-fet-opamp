magic
tech sky130A
magscale 1 2
timestamp 1712676954
<< metal3 >>
rect -1941 1512 1941 1540
rect -1941 -1512 1857 1512
rect 1921 -1512 1941 1512
rect -1941 -1540 1941 -1512
<< via3 >>
rect 1857 -1512 1921 1512
<< mimcap >>
rect -1901 1460 1609 1500
rect -1901 -1460 -1861 1460
rect 1569 -1460 1609 1460
rect -1901 -1500 1609 -1460
<< mimcapcontact >>
rect -1861 -1460 1569 1460
<< metal4 >>
rect 1841 1512 1937 1528
rect -1862 1460 1570 1461
rect -1862 -1460 -1861 1460
rect 1569 -1460 1570 1460
rect -1862 -1461 1570 -1460
rect 1841 -1512 1857 1512
rect 1921 -1512 1937 1512
rect 1841 -1528 1937 -1512
<< properties >>
string FIXED_BBOX -1941 -1540 1649 1540
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 17.55 l 15 val 538.869 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
