magic
tech sky130A
magscale 1 2
timestamp 1712682590
<< pwell >>
rect -468 -1372 32 -1262
<< locali >>
rect -1652 -136 -1470 -122
rect -1652 -192 -1638 -136
rect -1482 -192 -1470 -136
rect -1652 -982 -1470 -192
rect -1652 -1008 -1028 -982
rect -1650 -1038 -1028 -1008
rect -1650 -1260 -1470 -1038
rect -1650 -1380 -1614 -1260
rect -1504 -1380 -1470 -1260
rect -1650 -1420 -1470 -1380
<< viali >>
rect -418 140 -14 174
rect 1134 140 1520 174
rect -1206 30 -1042 66
rect 3250 10 3726 44
rect -1638 -192 -1482 -136
rect -420 -642 -14 -608
rect 1264 -642 1440 -608
rect -1614 -1380 -1504 -1260
rect 2394 -1358 2488 -1324
rect -356 -1564 -46 -1530
rect 1250 -1564 1460 -1530
rect 3224 -1822 3736 -1788
rect -1216 -2084 -1042 -2050
<< metal1 >>
rect -1230 410 -1030 600
rect -1230 312 -1028 410
rect 374 312 772 314
rect -1230 310 3178 312
rect -1230 224 3844 310
rect -1230 66 -1028 224
rect -1230 30 -1206 66
rect -1042 30 -1028 66
rect -1230 18 -1028 30
rect -782 174 404 224
rect -782 140 -418 174
rect -14 140 404 174
rect -782 20 404 140
rect 746 216 1940 224
rect 746 174 1938 216
rect 746 140 1134 174
rect 1520 140 1938 174
rect 746 20 1938 140
rect 2240 -14 2356 -6
rect 2240 -20 2248 -14
rect 1982 -22 2248 -20
rect -1392 -28 2248 -22
rect -1392 -80 -1384 -28
rect -1304 -64 2248 -28
rect -1304 -80 -1298 -64
rect -1392 -88 -1298 -80
rect 2240 -72 2248 -64
rect 2348 -72 2356 -14
rect 2240 -82 2356 -72
rect -1652 -136 -1470 -122
rect -1652 -192 -1638 -136
rect -1482 -152 -1470 -136
rect -788 -152 400 -114
rect -1482 -184 400 -152
rect -1482 -192 -1470 -184
rect -1652 -208 -1470 -192
rect -2332 -352 -2132 -284
rect -2332 -356 1000 -352
rect -2332 -416 860 -356
rect 992 -416 1000 -356
rect -2332 -420 1000 -416
rect -2332 -484 -2132 -420
rect 1234 -508 1478 -118
rect 1946 -360 2028 -352
rect 1946 -414 1954 -360
rect 2022 -414 2028 -360
rect 1946 -420 2028 -414
rect -468 -572 1478 -508
rect -468 -608 28 -572
rect -468 -642 -420 -608
rect -14 -642 28 -608
rect -2328 -790 -2128 -722
rect -468 -758 28 -642
rect 1234 -608 1478 -572
rect 1234 -642 1264 -608
rect 1440 -642 1478 -608
rect 1234 -754 1478 -642
rect -2328 -864 492 -790
rect 1988 -810 2028 -420
rect 662 -852 2028 -810
rect -2328 -922 -2128 -864
rect -868 -866 492 -864
rect 1988 -888 2028 -852
rect -2330 -1288 -2130 -1220
rect -1654 -1260 -1470 -1220
rect -1654 -1288 -1614 -1260
rect -2330 -1352 -1614 -1288
rect -2330 -1420 -2130 -1352
rect -1654 -1380 -1614 -1352
rect -1504 -1380 -1470 -1260
rect -468 -1324 32 -900
rect 1232 -1048 1480 -902
rect 1232 -1122 2372 -1048
rect 1232 -1272 1480 -1122
rect -858 -1374 2000 -1324
rect -1654 -1420 -1470 -1380
rect -468 -1530 32 -1414
rect -468 -1564 -356 -1530
rect -46 -1564 32 -1530
rect -1392 -2026 -1298 -2018
rect -1392 -2090 -1384 -2026
rect -1304 -2038 -1298 -2026
rect -1304 -2040 -1030 -2038
rect -468 -2040 32 -1564
rect 1230 -1530 1480 -1416
rect 1230 -1564 1250 -1530
rect 1460 -1564 1480 -1530
rect 1230 -2040 1480 -1564
rect 2138 -1558 2186 -1122
rect 2418 -1258 2474 224
rect 3148 44 3844 224
rect 3148 10 3250 44
rect 3726 10 3844 44
rect 2550 -18 2648 -8
rect 2550 -72 2558 -18
rect 2642 -72 2648 -18
rect 2550 -82 2648 -72
rect 2576 -154 2612 -82
rect 3148 -104 3844 10
rect 2576 -200 4188 -154
rect 3316 -796 3718 -248
rect 5420 -796 5620 -750
rect 3316 -908 5620 -796
rect 2508 -1020 2554 -1018
rect 2508 -1032 3094 -1020
rect 2508 -1138 2864 -1032
rect 3082 -1138 3094 -1032
rect 2508 -1154 3094 -1138
rect 2382 -1324 2512 -1316
rect 2382 -1358 2394 -1324
rect 2488 -1358 2512 -1324
rect 2382 -1368 2512 -1358
rect 2138 -1568 2224 -1558
rect 2138 -1628 2148 -1568
rect 2216 -1628 2224 -1568
rect 2138 -1638 2224 -1628
rect 2382 -2038 2510 -1368
rect 3316 -1530 3718 -908
rect 2564 -1564 2672 -1552
rect 2564 -1624 2574 -1564
rect 2660 -1574 2672 -1564
rect 2660 -1576 2876 -1574
rect 2660 -1618 4170 -1576
rect 2660 -1624 2672 -1618
rect 2564 -1636 2672 -1624
rect 3132 -1788 3834 -1674
rect 3132 -1822 3224 -1788
rect 3736 -1822 3834 -1788
rect 3132 -2038 3834 -1822
rect 4970 -1676 5174 -908
rect 5420 -950 5620 -908
rect 4970 -2004 4988 -1676
rect 5160 -2004 5174 -1676
rect 4970 -2022 5174 -2004
rect 2382 -2040 3834 -2038
rect -1304 -2050 3834 -2040
rect -1304 -2084 -1216 -2050
rect -1042 -2084 3834 -2050
rect -1304 -2090 3834 -2084
rect -1392 -2096 3834 -2090
rect -1392 -2098 3138 -2096
rect -1392 -2100 -1030 -2098
rect 2438 -2100 3138 -2098
rect -1230 -2552 -1030 -2100
<< via1 >>
rect -1384 -80 -1304 -28
rect 2248 -72 2348 -14
rect 860 -416 992 -356
rect 1954 -414 2022 -360
rect -1384 -2090 -1304 -2026
rect 2558 -72 2642 -18
rect 2864 -1138 3082 -1032
rect 2148 -1628 2216 -1568
rect 2574 -1624 2660 -1564
rect 4988 -2004 5160 -1676
<< metal2 >>
rect 2240 -14 2356 -6
rect -1392 -28 -1298 -22
rect -1392 -80 -1384 -28
rect -1304 -80 -1298 -28
rect -1392 -2026 -1298 -80
rect 2240 -72 2248 -14
rect 2348 -20 2356 -14
rect 2550 -18 2648 -8
rect 2550 -20 2558 -18
rect 2348 -64 2558 -20
rect 2348 -72 2356 -64
rect 2240 -82 2356 -72
rect 2550 -72 2558 -64
rect 2642 -72 2648 -18
rect 2550 -82 2648 -72
rect 846 -356 2028 -352
rect 846 -416 860 -356
rect 992 -360 2028 -356
rect 992 -414 1954 -360
rect 2022 -414 2028 -360
rect 992 -416 2028 -414
rect 846 -420 2028 -416
rect 2848 -1032 3094 -1020
rect 2848 -1138 2864 -1032
rect 3082 -1138 3094 -1032
rect 2848 -1154 3094 -1138
rect 2138 -1568 2224 -1558
rect 2138 -1628 2148 -1568
rect 2216 -1574 2224 -1568
rect 2564 -1564 2672 -1552
rect 2564 -1574 2574 -1564
rect 2216 -1620 2574 -1574
rect 2216 -1628 2224 -1620
rect 2138 -1638 2224 -1628
rect 2564 -1624 2574 -1620
rect 2660 -1624 2672 -1564
rect 2564 -1636 2672 -1624
rect 4970 -1676 5178 -1654
rect 4970 -2004 4988 -1676
rect 5160 -2004 5178 -1676
rect 4970 -2022 5178 -2004
rect -1392 -2090 -1384 -2026
rect -1304 -2090 -1298 -2026
rect -1392 -2100 -1298 -2090
<< via2 >>
rect 2864 -1138 3082 -1032
rect 4988 -2004 5160 -1676
<< metal3 >>
rect 2848 -1032 3094 -1020
rect 2848 -1138 2864 -1032
rect 3082 -1138 3094 -1032
rect 2848 -1154 3094 -1138
rect 4970 -1676 5178 -1654
rect 4970 -2004 4988 -1676
rect 5160 -2004 5178 -1676
rect 4970 -2022 5178 -2004
<< via3 >>
rect 2864 -1138 3082 -1032
rect 4988 -2004 5160 -1676
<< metal4 >>
rect 4490 -1022 4622 -1020
rect 2848 -1032 4622 -1022
rect 2848 -1138 2864 -1032
rect 3082 -1138 4622 -1032
rect 2848 -1156 4622 -1138
rect 4490 -2402 4622 -1156
rect 2704 -2474 4622 -2402
rect 4974 -1676 5176 -1656
rect 4974 -2004 4988 -1676
rect 5160 -2004 5176 -1676
rect 2704 -3796 2764 -2474
rect 4974 -2758 5176 -2004
rect 2704 -3874 3066 -3796
use sky130_fd_pr__res_generic_l1_SQKU9V  R1
timestamp 1712505088
transform 1 0 -1128 0 1 -481
box -100 -557 100 557
use sky130_fd_pr__res_generic_l1_SQKU9V  R2
timestamp 1712505088
transform 1 0 -1128 0 1 -1539
box -100 -557 100 557
use sky130_fd_pr__cap_mim_m3_1_QJVKAD  sky130_fd_pr__cap_mim_m3_1_QJVKAD_0
timestamp 1712676954
transform 0 -1 4520 1 0 -4679
box -1941 -1540 1941 1540
use sky130_fd_pr__pfet_01v8_XPP7BA  XM1
timestamp 1712505088
transform 0 1 -189 -1 0 -828
box -256 -819 256 819
use sky130_fd_pr__pfet_01v8_XPP7BA  XM2
timestamp 1712505088
transform 0 1 1343 -1 0 -828
box -256 -819 256 819
use sky130_fd_pr__nfet_01v8_3BHWKV  XM3
timestamp 1712505088
transform 0 1 -186 -1 0 -1344
box -256 -810 256 810
use sky130_fd_pr__nfet_01v8_3BHWKV  XM4
timestamp 1712505088
transform 0 1 1328 -1 0 -1344
box -256 -810 256 810
use sky130_fd_pr__pfet_01v8_XPP7BA  XM5
timestamp 1712505088
transform 0 1 1343 -1 0 -46
box -256 -819 256 819
use sky130_fd_pr__nfet_01v8_3BHWKV  XM6
timestamp 1712505088
transform 0 1 3500 -1 0 -1602
box -256 -810 256 810
use sky130_fd_pr__pfet_01v8_XPP7BA  XM7
timestamp 1712505088
transform 0 1 3509 -1 0 -176
box -256 -819 256 819
use sky130_fd_pr__pfet_01v8_XPP7BA  XM8
timestamp 1712505088
transform 0 1 -189 -1 0 -46
box -256 -819 256 819
use sky130_fd_pr__nfet_01v8_7QHW3M  XM9
timestamp 1712505088
transform 1 0 2442 0 1 -1084
box -256 -310 256 310
<< labels >>
flabel metal1 -1230 400 -1030 600 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 -2330 -1420 -2130 -1220 0 FreeSans 256 0 0 0 ZREF
port 1 nsew
flabel metal1 -1230 -2552 -1030 -2352 0 FreeSans 256 0 0 0 VGND
port 5 nsew
flabel metal1 -2328 -922 -2128 -722 0 FreeSans 256 0 0 0 vin_n
port 2 nsew
flabel metal1 -2332 -484 -2132 -284 0 FreeSans 256 0 0 0 vin_p
port 3 nsew
flabel metal1 5420 -950 5620 -750 0 FreeSans 256 0 0 0 Vout
port 4 nsew
<< end >>
