magic
tech sky130A
timestamp 1712505088
<< pwell >>
rect -128 -155 128 155
<< nmos >>
rect -30 -50 30 50
<< ndiff >>
rect -59 44 -30 50
rect -59 -44 -53 44
rect -36 -44 -30 44
rect -59 -50 -30 -44
rect 30 44 59 50
rect 30 -44 36 44
rect 53 -44 59 44
rect 30 -50 59 -44
<< ndiffc >>
rect -53 -44 -36 44
rect 36 -44 53 44
<< psubdiff >>
rect -110 120 -62 137
rect 62 120 110 137
rect -110 89 -93 120
rect 93 89 110 120
rect -110 -120 -93 -89
rect 93 -120 110 -89
rect -110 -137 -62 -120
rect 62 -137 110 -120
<< psubdiffcont >>
rect -62 120 62 137
rect -110 -89 -93 89
rect 93 -89 110 89
rect -62 -137 62 -120
<< poly >>
rect -30 86 30 94
rect -30 69 -22 86
rect 22 69 30 86
rect -30 50 30 69
rect -30 -69 30 -50
rect -30 -86 -22 -69
rect 22 -86 30 -69
rect -30 -94 30 -86
<< polycont >>
rect -22 69 22 86
rect -22 -86 22 -69
<< locali >>
rect -110 120 -62 137
rect 62 120 110 137
rect -110 89 -93 120
rect 93 89 110 120
rect -30 69 -22 86
rect 22 69 30 86
rect -53 44 -36 52
rect -53 -52 -36 -44
rect 36 44 53 52
rect 36 -52 53 -44
rect -30 -86 -22 -69
rect 22 -86 30 -69
rect -110 -120 -93 -89
rect 93 -120 110 -89
rect -110 -137 -62 -120
rect 62 -137 110 -120
<< viali >>
rect -22 69 22 86
rect -53 -44 -36 44
rect 36 -44 53 44
rect -22 -86 22 -69
<< metal1 >>
rect -28 86 28 89
rect -28 69 -22 86
rect 22 69 28 86
rect -28 66 28 69
rect -56 44 -33 50
rect -56 -44 -53 44
rect -36 -44 -33 44
rect -56 -50 -33 -44
rect 33 44 56 50
rect 33 -44 36 44
rect 53 -44 56 44
rect 33 -50 56 -44
rect -28 -69 28 -66
rect -28 -86 -22 -69
rect 22 -86 28 -69
rect -28 -89 28 -86
<< properties >>
string FIXED_BBOX -101 -128 101 128
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 0.6 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
