** sch_path: /home/dsatizabal/tt06-fet-opamp/xschem/opamp_tb.sch
**.subckt opamp_tb
x1 net2 GND net1 Vi Vo net3 opamp
R1 net1 GND 1k m=1
R2 Vo net1 2k m=1
V1 Vi GND sin(0 20m 100) ac 1
V3 net2 net3 1.8
x1 net5 GND net4 Vilay Volay net6 opamp_parax
R3 net4 GND 1k m=1
R4 Volay net4 2k m=1
V2 Vilay GND sin(0 20m 100) ac 1
V4 net5 net6 1.8
**** begin user architecture code



.control
tran 10u 100m
write opamp_tb.raw
ac dec 100 1 100MEG
write opamp_tb_ac.raw
.endc




.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/dsatizabal/zerotoasic/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/dsatizabal/zerotoasic/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/dsatizabal/zerotoasic/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/dsatizabal/zerotoasic/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends

* expanding   symbol:  opamp.sym # of pins=6
** sym_path: /home/dsatizabal/tt06-fet-opamp/xschem/opamp.sym
** sch_path: /home/dsatizabal/tt06-fet-opamp/xschem/opamp.sch
.subckt opamp VDD ZREF vin_n vin_p Vout VGND
*.ipin vin_n
*.ipin vin_p
*.opin Vout
*.iopin VDD
*.iopin ZREF
*.iopin VGND
XM1 net1 vin_n net3 net3 sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net2 vin_p net3 net3 sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net1 net1 VGND VGND sky130_fd_pr__nfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net2 net1 VGND VGND sky130_fd_pr__nfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net3 VGND VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 Vout VGND VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 ZREF VGND VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 net4 VDD net2 VGND sky130_fd_pr__nfet_01v8 L=0.6 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC1 net4 Vout sky130_fd_pr__cap_mim_m3_1 W=17.55 L=15 MF=6 m=6
XM6 Vout net2 VGND VGND sky130_fd_pr__nfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
R1 ZREF VDD sky130_fd_pr__res_generic_l1 W=1 L=5 m=1
R2 VGND ZREF sky130_fd_pr__res_generic_l1 W=1 L=5 m=1
.ends


* expanding   symbol:  opamp_parax.sym # of pins=6
** sym_path: /home/dsatizabal/tt06-fet-opamp/xschem/opamp.sym
.include /home/dsatizabal/tt06-fet-opamp/mag/opamp.sim.spice
.GLOBAL GND
.end
