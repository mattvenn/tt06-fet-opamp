magic
tech sky130A
timestamp 1712505088
<< pwell >>
rect -128 -405 128 405
<< nmos >>
rect -30 -300 30 300
<< ndiff >>
rect -59 294 -30 300
rect -59 -294 -53 294
rect -36 -294 -30 294
rect -59 -300 -30 -294
rect 30 294 59 300
rect 30 -294 36 294
rect 53 -294 59 294
rect 30 -300 59 -294
<< ndiffc >>
rect -53 -294 -36 294
rect 36 -294 53 294
<< psubdiff >>
rect -110 370 -62 387
rect 62 370 110 387
rect -110 339 -93 370
rect 93 339 110 370
rect -110 -370 -93 -339
rect 93 -370 110 -339
rect -110 -387 -62 -370
rect 62 -387 110 -370
<< psubdiffcont >>
rect -62 370 62 387
rect -110 -339 -93 339
rect 93 -339 110 339
rect -62 -387 62 -370
<< poly >>
rect -30 336 30 344
rect -30 319 -22 336
rect 22 319 30 336
rect -30 300 30 319
rect -30 -319 30 -300
rect -30 -336 -22 -319
rect 22 -336 30 -319
rect -30 -344 30 -336
<< polycont >>
rect -22 319 22 336
rect -22 -336 22 -319
<< locali >>
rect -110 370 -62 387
rect 62 370 110 387
rect -110 339 -93 370
rect 93 339 110 370
rect -30 319 -22 336
rect 22 319 30 336
rect -53 294 -36 302
rect -53 -302 -36 -294
rect 36 294 53 302
rect 36 -302 53 -294
rect -30 -336 -22 -319
rect 22 -336 30 -319
rect -110 -370 -93 -339
rect 93 -370 110 -339
rect -110 -387 -62 -370
rect 62 -387 110 -370
<< viali >>
rect -22 319 22 336
rect -53 -294 -36 294
rect 36 -294 53 294
rect -22 -336 22 -319
<< metal1 >>
rect -28 336 28 339
rect -28 319 -22 336
rect 22 319 28 336
rect -28 316 28 319
rect -56 294 -33 300
rect -56 -294 -53 294
rect -36 -294 -33 294
rect -56 -300 -33 -294
rect 33 294 56 300
rect 33 -294 36 294
rect 53 -294 56 294
rect 33 -300 56 -294
rect -28 -319 28 -316
rect -28 -336 -22 -319
rect 22 -336 28 -319
rect -28 -339 28 -336
<< properties >>
string FIXED_BBOX -101 -378 101 378
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 6.0 l 0.6 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
