magic
tech sky130A
magscale 1 2
timestamp 1712505088
<< metal3 >>
rect -1941 9812 1941 9840
rect -1941 6788 1857 9812
rect 1921 6788 1941 9812
rect -1941 6760 1941 6788
rect -1941 6492 1941 6520
rect -1941 3468 1857 6492
rect 1921 3468 1941 6492
rect -1941 3440 1941 3468
rect -1941 3172 1941 3200
rect -1941 148 1857 3172
rect 1921 148 1941 3172
rect -1941 120 1941 148
rect -1941 -148 1941 -120
rect -1941 -3172 1857 -148
rect 1921 -3172 1941 -148
rect -1941 -3200 1941 -3172
rect -1941 -3468 1941 -3440
rect -1941 -6492 1857 -3468
rect 1921 -6492 1941 -3468
rect -1941 -6520 1941 -6492
rect -1941 -6788 1941 -6760
rect -1941 -9812 1857 -6788
rect 1921 -9812 1941 -6788
rect -1941 -9840 1941 -9812
<< via3 >>
rect 1857 6788 1921 9812
rect 1857 3468 1921 6492
rect 1857 148 1921 3172
rect 1857 -3172 1921 -148
rect 1857 -6492 1921 -3468
rect 1857 -9812 1921 -6788
<< mimcap >>
rect -1901 9760 1609 9800
rect -1901 6840 -1861 9760
rect 1569 6840 1609 9760
rect -1901 6800 1609 6840
rect -1901 6440 1609 6480
rect -1901 3520 -1861 6440
rect 1569 3520 1609 6440
rect -1901 3480 1609 3520
rect -1901 3120 1609 3160
rect -1901 200 -1861 3120
rect 1569 200 1609 3120
rect -1901 160 1609 200
rect -1901 -200 1609 -160
rect -1901 -3120 -1861 -200
rect 1569 -3120 1609 -200
rect -1901 -3160 1609 -3120
rect -1901 -3520 1609 -3480
rect -1901 -6440 -1861 -3520
rect 1569 -6440 1609 -3520
rect -1901 -6480 1609 -6440
rect -1901 -6840 1609 -6800
rect -1901 -9760 -1861 -6840
rect 1569 -9760 1609 -6840
rect -1901 -9800 1609 -9760
<< mimcapcontact >>
rect -1861 6840 1569 9760
rect -1861 3520 1569 6440
rect -1861 200 1569 3120
rect -1861 -3120 1569 -200
rect -1861 -6440 1569 -3520
rect -1861 -9760 1569 -6840
<< metal4 >>
rect -198 9761 -94 9960
rect 1837 9812 1941 9960
rect -1862 9760 1570 9761
rect -1862 6840 -1861 9760
rect 1569 6840 1570 9760
rect -1862 6839 1570 6840
rect -198 6441 -94 6839
rect 1837 6788 1857 9812
rect 1921 6788 1941 9812
rect 1837 6492 1941 6788
rect -1862 6440 1570 6441
rect -1862 3520 -1861 6440
rect 1569 3520 1570 6440
rect -1862 3519 1570 3520
rect -198 3121 -94 3519
rect 1837 3468 1857 6492
rect 1921 3468 1941 6492
rect 1837 3172 1941 3468
rect -1862 3120 1570 3121
rect -1862 200 -1861 3120
rect 1569 200 1570 3120
rect -1862 199 1570 200
rect -198 -199 -94 199
rect 1837 148 1857 3172
rect 1921 148 1941 3172
rect 1837 -148 1941 148
rect -1862 -200 1570 -199
rect -1862 -3120 -1861 -200
rect 1569 -3120 1570 -200
rect -1862 -3121 1570 -3120
rect -198 -3519 -94 -3121
rect 1837 -3172 1857 -148
rect 1921 -3172 1941 -148
rect 1837 -3468 1941 -3172
rect -1862 -3520 1570 -3519
rect -1862 -6440 -1861 -3520
rect 1569 -6440 1570 -3520
rect -1862 -6441 1570 -6440
rect -198 -6839 -94 -6441
rect 1837 -6492 1857 -3468
rect 1921 -6492 1941 -3468
rect 1837 -6788 1941 -6492
rect -1862 -6840 1570 -6839
rect -1862 -9760 -1861 -6840
rect 1569 -9760 1570 -6840
rect -1862 -9761 1570 -9760
rect -198 -9960 -94 -9761
rect 1837 -9812 1857 -6788
rect 1921 -9812 1941 -6788
rect 1837 -9960 1941 -9812
<< properties >>
string FIXED_BBOX -1941 6760 1649 9840
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 17.55 l 15.0 val 538.869 carea 2.00 cperi 0.19 nx 1 ny 6 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
